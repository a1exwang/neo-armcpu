/*
 * $File: int_def.vh
 * $Date: Fri Dec 20 11:36:21 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

// definition of interrupt numbers

`define INT_TIMER	7
`define INT_KBD		6
`define INT_SL811   5
`define INT_COM		4

// vim: ft=verilog


